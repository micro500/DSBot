--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   20:16:55 08/06/2015
-- Design Name:   
-- Module Name:   E:/FPGA/DS_Bot/main_test.vhd
-- Project Name:  DS_Bot
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: main
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY main_test IS
END main_test;
 
ARCHITECTURE behavior OF main_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT main
    PORT(
         clk : IN  std_logic;
         sclk : IN  std_logic;
         en : IN  std_logic;
         di : IN  std_logic;
         do : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal sclk : std_logic := '1';
   signal en : std_logic := '1';
   signal di : std_logic := '1';

 	--Outputs
   signal do : std_logic;

   -- Clock period definitions
   constant clk_period : time := 32.25 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: main PORT MAP (
          clk => clk,
          sclk => sclk,
          en => en,
          di => di,
          do => do
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
      
      
wait for 1000ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 600ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 750ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '1';
di <= '1';
wait for 16749475ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 25ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 575ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 725ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '1';
di <= '1';
wait for 16658400ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 575ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 750ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '1';
di <= '1';
wait for 16706875ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '1';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '1';
wait for 25ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 600ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 750ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '0';
en <= '0';
di <= '0';
wait for 225ns;
sclk <= '1';
en <= '0';
di <= '0';
wait for 250ns;
sclk <= '1';
en <= '1';
di <= '1';






      wait;
   end process;

END;
